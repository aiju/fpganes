`timescale 1 ns / 1 ps
`default_nettype none

`define VRAMINC 2
`define SPRTAB 3
`define PATTAB 4
`define SPR16 5
`define GENNMI 7

`define GRAY 0
`define BG8 1
`define SPR8 2
`define SHOWBG 3
`define SHOWSPR 4
`define INTR 5
`define INTG 6
`define INTB 7

`define MIRRHOR 0
`define MIRRVER 1
`define MIRRA 2
`define MIRRB 3
`define MIRR4 4
