`include "dat.vh"

module tickgen(
	input wire clk,
	input wire stall,
	output reg cputick,
	output reg pputick
);

	

endmodule
